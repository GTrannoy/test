--_________________________________________________________________________________________________
--                                                                                                |
--                                        |The nanoFIP|                                           |
--                                                                                                |
--                                        CERN,BE/CO-HT                                           |
--________________________________________________________________________________________________|
--________________________________________________________________________________________________|

---------------------------------------------------------------------------------------------------
--! @file WF_manch_encoder.vhd                                                                    |
---------------------------------------------------------------------------------------------------

--! standard library
library IEEE; 

--! standard packages
use IEEE.STD_LOGIC_1164.all;  --! std_logic definitions
use IEEE.NUMERIC_STD.all;     --! conversion functions

---------------------------------------------------------------------------------------------------
--                                                                                               --
--                                       WF_manch_encoder                                        --
--                                                                                               --
---------------------------------------------------------------------------------------------------
--
--
--! @brief     Encoding of a word to its Manchester 2 (manch.) equivalent.
--!            This code ensures that there is one transition for each bit.
--!            bit            :    "0"           "1"
--!            manch. encoded :   "0 1"         "1 0"
--!            scheme         :    _|-           -|_
--
--
--! @author    Pablo Alvarez Sanchez (Pablo.Alvarez.Sanchez@cern.ch)\n
--!            Evangelia Gousiou     (Evangelia.Gousiou@cern.ch)    \n
--
--
--! @date      10/12/2010
--
--
--! @version   v0.02
--
--
--! @details \n  
--
--!   \n<b>Dependencies:</b>\n
--
--
--!   \n<b>Modified by:</b>   \n
--!     Evangelia Gousiou     \n
--
--------------------------------------------------------------------------------------------------- 
--
--!   \n\n<b>Last changes:</b>\n
--!     -> 11/2010  v0.01  EG  1st version           \n
--!     -> 12/2010  v0.02  EG  cleaned-up, commented \n
--! 
--
--------------------------------------------------------------------------------------------------- 
--
--! @todo 
--!   -> 
--
--------------------------------------------------------------------------------------------------- 

---/!\----------------------------/!\----------------------------/!\-------------------------/!\---
--                               Synplify Premier D-2009.12 Warnings                             --
-- -- --  --  --  --  --  --  --  --  --  --  --  --  --  --  -- --  --  --  --  --  --  --  --  --
--                                         No Warnings                                           --
---------------------------------------------------------------------------------------------------


--=================================================================================================
--!                           Entity declaration for WF_manch_encoder
--=================================================================================================

entity WF_manch_encoder is

  generic (word_length : natural := 8);                               --! default word length: 8
  port (
  -- INPUT 
    word_i       : in  std_logic_vector(word_length-1 downto 0);      --! input word        


  -- OUTPUT
    word_manch_o : out std_logic_vector((2*word_length)-1 downto 0)   --! output encoded word
      );
end entity WF_manch_encoder;


--=================================================================================================
--!                                  architecture declaration
--=================================================================================================
architecture rtl of WF_manch_encoder is


--=================================================================================================
--                                       architecture begin
--=================================================================================================  
begin

---------------------------------------------------------------------------------------------------
--! @brief Combinatorial process Manchester_Encoder: The process takes a word (ex. 8 bits) and
--! creates its manchester encoded equivalent (ex. 16 bits).
--! Each bit '1' is replaced by '10' and each bit '0' by '01'. 

  Manchester_Encoder: process (word_i)
  begin

    for I in word_i'range loop

      word_manch_o(I*2)   <= not word_i(I);

      word_manch_o(I*2+1) <= word_i(I);

    end loop;
  end process;


end architecture rtl;
--=================================================================================================
--                                      architecture end
--=================================================================================================
---------------------------------------------------------------------------------------------------
--                                    E N D   O F   F I L E
---------------------------------------------------------------------------------------------------